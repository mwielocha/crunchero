create keyspace ProfileService
with placement_strategy = 'org.apache.cassandra.locator.NetworkTopologyStrategy'
and strategy_options={datacenter1:3};

